`timescale  1ns / 1ps

module tb_stream_demux;

// stream_demux Parameters
parameter PERIOD   = 10;
parameter DATA_WD  = 32;

// stream_demux Inputs
reg   clk                   ;
reg   rstn                  ;
reg   sel                   ;
reg   [DATA_WD-1:0]  a_data ;
reg   a_valid               ;
reg   b_ready               ;
reg   c_ready               ;

// stream_demux Outputs
wire  a_ready                              ;
wire  [DATA_WD-1:0]  b_data                ;
wire  b_valid                              ;
wire  [DATA_WD-1:0]  c_data                ;
wire  c_valid                              ;

//fire 
wire  a_fire,b_fire,c_fire;
assign a_fire = a_valid && a_ready;
assign b_fire = b_valid && b_ready;
assign c_fire = c_valid && c_ready;


initial
begin
    clk = 0;
    forever #(PERIOD/2)  clk=~clk;
end

initial
begin
    rstn = 0;
    #(PERIOD*2) rstn  =  1;
end


initial begin
    $dumpfile("test.vcd");
    $dumpvars;
end

always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        a_valid <= 1'b0;
        a_data <= 'b0;
        //b_valid <= 1'b0;
        //b_data <= 'b0;
        sel <= 1'b0;   
    end
    else begin
        /*if (!a_valid) begin
            a_valid <= $random;
        end
        else if (a_valid && a_ready) begin
            a_valid <= $random;
            a_data <= a_data + 1'b1;           
        end*/
        if (!a_valid || a_ready) begin
            a_valid <= $random;
            if (a_valid) begin
                a_data <= a_data + 1;
            end
        end
        sel <= sel + a_fire;

    end
end

always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        c_ready <= 1'b1;
        b_ready <= 1'b1;
    end
    else begin
        b_ready <= $random;
        c_ready <= $random;
    end
end


stream_demux #(
    .DATA_WD ( DATA_WD ))
 u_stream_demux (
    .clk                     ( clk                    ),
    .rstn                    ( rstn                   ),
    .sel                     ( sel                    ),
    .a_data                  ( a_data   [DATA_WD-1:0] ),
    .a_valid                 ( a_valid                ),
    .b_ready                 ( b_ready                ),
    .c_ready                 ( c_ready                ),

    .a_ready                 ( a_ready                ),
    .b_data                  ( b_data   [DATA_WD-1:0] ),
    .b_valid                 ( b_valid                ),
    .c_data                  ( c_data   [DATA_WD-1:0] ),
    .c_valid                 ( c_valid                )
);

initial
begin
    #5000;
    $finish;
end

endmodule